`timescale 1ns / 1ps
module Pipelined_MIPS32(clk1 ,clk2);
input clk1,clk2;
reg [31:0] PC,IF_ID_IR,IF_ID_NPC; //btw IF,ID
reg [31:0] ID_EX_IR,ID_EX_NPC,ID_EX_A,ID_EX_B,ID_EX_Imm; //btw ID,EX
reg [31:0] EX_MEM_IR,EX_MEM_B,EX_MEM_ALUOUT; //btw EX,MEM
reg EX_MEM_cond;
reg [31:0] MEM_WB_ALUOUT,MEM_WB_IR,MEM_WB_LMD; //btw MEM,WB
reg [2:0] ID_EX_TYPE ,EX_MEM_TYPE,MEM_WB_TYPE; //for type of instruction
reg [31:0] regbank[0:31];
reg [31:0] instr_mem[0:1023]; // Instruction memory
reg [31:0] data_mem[0:1023];  // Data memory
parameter ADD=  6'b000000,
          SUB=  6'b000001,
          AND=  6'b000010,
          OR=   6'b000011,
          SLT=  6'b000100,
          MUL=  6'b000101,
          HLT=  6'b111111,
          LW=   6'b001000,
          SW=   6'b001001,
          ADDI= 6'b001010,
          SUBI= 6'b001011,
          SLTI= 6'b001100,
          BNEQZ=6'b001101,
          BEQZ= 6'b001110;  
parameter RR_ALU=3'b000,
          RM_ALU=3'b001,
          LOAD=3'b010,
          STORE=3'b011,
          BRANCH=3'b100,
          HALT=3'b101;
reg HALTED;
reg TAKEN_BRANCH;
initial begin
          PC = 0;
          HALTED = 0;
          TAKEN_BRANCH = 0;
end
//IF STAGE 
always@(posedge clk1)
    if(!HALTED)
    begin
        if(((EX_MEM_IR[31:26]==BEQZ)&&(EX_MEM_cond==1)) || ((EX_MEM_IR[31:26]==BNEQZ)&&(EX_MEM_cond==0)))
            begin
                IF_ID_IR    <=instr_mem[EX_MEM_ALUOUT];
                TAKEN_BRANCH<=1'b1;
                IF_ID_NPC   <=EX_MEM_ALUOUT+1;
                PC          <=EX_MEM_ALUOUT+1;
            end
        else
            begin
                IF_ID_IR <=instr_mem[PC];
                IF_ID_NPC<=PC+1;
                PC       <=PC+1;
            end
    end
//ID STAGE 
always@(posedge clk2)
    if(HALTED==0)
    begin 
        if (IF_ID_IR[25:21]==5'b00000)
                ID_EX_A<=0;
        else
                ID_EX_A<=regbank[IF_ID_IR[25:21]];
        if (IF_ID_IR[20:16]==5'b00000)
                ID_EX_B<=0;
        else
                ID_EX_B<=regbank[IF_ID_IR[20:16]];    
                
     ID_EX_NPC<=IF_ID_NPC;
     ID_EX_IR<=IF_ID_IR;
     ID_EX_Imm<={{16{IF_ID_IR[15]}},{IF_ID_IR[15:0]}};
     case(IF_ID_IR[31:26]) //to identify type of operation
       ADD,SUB,MUL,AND,OR,SLT : ID_EX_TYPE<= RR_ALU;
       ADDI,SUBI,SLTI:          ID_EX_TYPE<= RM_ALU; 
       LW:                      ID_EX_TYPE<=LOAD;
       SW:                      ID_EX_TYPE<=STORE;
       BNEQZ,BEQZ:              ID_EX_TYPE<=BRANCH;
       HLT:                     ID_EX_TYPE<=HALT;
       default:                 ID_EX_TYPE<=HALT;
     endcase
    end
//EX STAGE
always@(posedge clk1)
begin
  if(!HALTED)
  begin
    EX_MEM_TYPE<=ID_EX_TYPE;
    EX_MEM_IR<=ID_EX_IR;
    TAKEN_BRANCH<=0;
    
    case(ID_EX_TYPE)
    RR_ALU : begin
               case(ID_EX_IR[31:26])
                    ADD : EX_MEM_ALUOUT <= ID_EX_A+ID_EX_B;
                    SUB : EX_MEM_ALUOUT <= ID_EX_A-ID_EX_B;
                    MUL : EX_MEM_ALUOUT <= ID_EX_A*ID_EX_B;
                    AND : EX_MEM_ALUOUT <=ID_EX_A & ID_EX_B;
                    OR : EX_MEM_ALUOUT <= ID_EX_A | ID_EX_B;
                    SLT : EX_MEM_ALUOUT <=(ID_EX_A < ID_EX_B)? 32'd1 : 32'd0;
                    default : EX_MEM_ALUOUT <=32'hxxxxxxxx;
                endcase
             end
    RM_ALU : begin
               case(ID_EX_IR[31:26])
                    ADDI: EX_MEM_ALUOUT<=ID_EX_A + ID_EX_Imm;
                    SUBI: EX_MEM_ALUOUT<=ID_EX_A - ID_EX_Imm;
                    SLTI:EX_MEM_ALUOUT <=(ID_EX_A < ID_EX_Imm)? 32'd1 : 32'd0;
                    default : EX_MEM_ALUOUT<= 32'hxxxxxxxx;
               endcase
             end
    LOAD ,STORE:
             begin
                    EX_MEM_ALUOUT<=ID_EX_A+ID_EX_Imm;
                    EX_MEM_B<=ID_EX_B;
             end
    BRANCH : begin
                   EX_MEM_cond<=(ID_EX_A==0);
                   EX_MEM_ALUOUT<=ID_EX_NPC+ID_EX_Imm;
             end
    endcase
  end
end
//MEM STAGE
always@(posedge clk2)
if(HALTED==0)
  begin
    MEM_WB_TYPE<=EX_MEM_TYPE;
    MEM_WB_IR<=EX_MEM_IR;
    case(EX_MEM_TYPE)
    RR_ALU,RM_ALU : 
                MEM_WB_ALUOUT<=EX_MEM_ALUOUT;
    LOAD :      MEM_WB_LMD<=data_mem[EX_MEM_ALUOUT];
    STORE:      if(TAKEN_BRANCH==0)
                   data_mem[EX_MEM_ALUOUT]<=EX_MEM_B;
    endcase
  end
//WB STAGE
always@(posedge clk1)
begin
  if(!TAKEN_BRANCH)
  case(MEM_WB_TYPE)
    RR_ALU : regbank[MEM_WB_IR[15:11]]<= MEM_WB_ALUOUT;
    RM_ALU : regbank[MEM_WB_IR[20:16]]<= MEM_WB_ALUOUT;
    LOAD   : regbank[MEM_WB_IR[20:16]]<= MEM_WB_LMD;
    HALT   : HALTED<=1'b1;
   endcase
end
endmodule

